--
-- VHDL Package Header RISCV_lib.ISA
--
-- Created:
--          by - flxbrggr.meyer (pc084)
--          at - 14:21:44 05/17/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
PACKAGE ISA IS
  ------------------------------------------
  -- ISA
  ------------------------------------------ 
  constant NOP: bit_vector :=b"00000" ;
END ISA;
