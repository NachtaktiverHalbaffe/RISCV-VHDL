--
-- VHDL Architecture RISCV_lib.mux_fw_rs2.behav
--
-- Created:
--          by - flxbrggr.meyer (pc084)
--          at - 14:58:26 05/31/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF mux_fw_rs2 IS
BEGIN
END ARCHITECTURE behav;

