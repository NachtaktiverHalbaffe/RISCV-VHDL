--
-- VHDL Architecture RISCV_lib.SdCardCtrl.behav
--
-- Created:
--          by - flxbrggr.meyer (pc084)
--          at - 17:19:50 07/12/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF SdCardCtrl IS
BEGIN
END ARCHITECTURE behav;

