--
-- VHDL Architecture RISCV_lib.Imm_Gen.behave
--
-- Created:
--          by - flxbrggr.meyer (pc085)
--          at - 17:54:55 05/10/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behave OF Imm_Gen IS
BEGIN
END ARCHITECTURE behave;

