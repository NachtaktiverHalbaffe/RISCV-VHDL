--
-- VHDL Architecture RISCV_lib.me_reg.behave
--
-- Created:
--          by - flxbrggr.meyer (pc085)
--          at - 17:55:36 05/10/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behave OF me_reg IS
BEGIN
END ARCHITECTURE behave;

