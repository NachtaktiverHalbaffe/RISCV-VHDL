--
-- VHDL Architecture RISCV_lib.mux_bpu_ra.behav
--
-- Created:
--          by - flxbrggr.meyer (pc084)
--          at - 10:53:36 06/28/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF mux_bpu_ra IS
BEGIN
END ARCHITECTURE behav;

