--
-- VHDL Entity RISCV_lib.WB_base.arch_name
--
-- Created:
--          by - flxbrggr.meyer (pc085)
--          at - 14:13:21 05/10/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity WB_base is
end entity WB_base;