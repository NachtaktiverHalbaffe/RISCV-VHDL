--
-- VHDL Architecture RISCV_lib.if_reg.behav
--
-- Created:
--          by - flxbrggr.meyer (pc085)
--          at - 17:52:35 05/10/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF if_reg IS
BEGIN
END ARCHITECTURE behav;

